module bitwise_not (
    B, data_result
);

    input [31:0] B;
    output [31:0] data_result;

    not Not0(data_result[0], B[0]);
    not Not1(data_result[1], B[1]);  
    not Not2(data_result[2], B[2]);  
    not Not3(data_result[3], B[3]);  
    not Not4(data_result[4], B[4]);  
    not Not5(data_result[5], B[5]);  
    not Not6(data_result[6], B[6]);  
    not Not7(data_result[7], B[7]);  
    not Not8(data_result[8], B[8]);  
    not Not9(data_result[9], B[9]);  
    not Not10(data_result[10], B[10]);  
    not Not11(data_result[11], B[11]);  
    not Not12(data_result[12], B[12]);  
    not Not13(data_result[13], B[13]);  
    not Not14(data_result[14], B[14]);  
    not Not15(data_result[15], B[15]);  
    not Not16(data_result[16], B[16]);  
    not Not17(data_result[17], B[17]);  
    not Not18(data_result[18], B[18]);  
    not Not19(data_result[19], B[19]);  
    not Not20(data_result[20], B[20]);  
    not Not21(data_result[21], B[21]);  
    not Not22(data_result[22], B[22]);  
    not Not23(data_result[23], B[23]);  
    not Not24(data_result[24], B[24]);  
    not Not25(data_result[25], B[25]);  
    not Not26(data_result[26], B[26]);  
    not Not27(data_result[27], B[27]);  
    not Not28(data_result[28], B[28]);  
    not Not29(data_result[29], B[29]);  
    not Not30(data_result[30], B[30]);  
    not Not31(data_result[31], B[31]);  

endmodule